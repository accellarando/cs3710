module cpuWithDatapath #(parameter size=16, NUMREGS=16)
	(input clk,
		reset, nextStateButton,
		output[9:0] leds,
		output[6:0] readData,
		output[6:0] writeData)
		
	stateMachine fsm(kjlkjlkjlkjlkjlkjjlkhojbihogugu80t70tgugjihjk);
endmodule 