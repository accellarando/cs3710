module datapath #(parameter SIZE = 16) (
	);