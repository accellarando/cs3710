`timescale 1ns / 1ps

module datapath_tb();
	/* Inputs */
//	reg 			clk, reset;
//	reg			writeEn;
//	reg[15:0] 	writeData;
//	reg[3:0] 	srcAddr, dstAddr;
//	integer 		counter;
//	
//	/* Outputs */
//	wire[15:0] 	readData1, readData2;
//	
//	/* Outputs */
//	/* Instantiate the Unit Under Test (UUT) */
//	registerFile uut (
//		.clk(clk),
//		.reset(reset),
//		.writeEn(writeEn),
//		.writeData(writeData),
//		.srcAddr(srcAddr),
//		.dstAddr(dstAddr),
//		.readData1(readData1),
//		.readData2(readData2)
//	);
	

endmodule
