module decoder 
	(
		input [4:0] flags_out,
		input [15:0] instr_out,
		output [4:0] rDest_in,
		output [15:0] alu_immed,
		output [7:0] opcodes,
		output [3:0] mux1_en, mux2_en,
		output [2:0] inst_type,
		output writeback_en
	)


endmodule

