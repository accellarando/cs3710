module stateMachine_tb();