module FSM
	(
		input clk, reset, writeback_en,
		input [1:0] inst_type,
		output addr_en, alu_mux_en, bus_mux_en, rDest_en, PC_en, mem_en, inst_en, flag_en, ram1_en, PC_count_en
	)
	
	

endmodule


// (clk, reset, writeback_en, inst_type, addr_en, alu_mux_en, bus_mux_en, rDest_en, PC_en, mem_en, inst_en, flag_en, ram1_en, PC_count_en);