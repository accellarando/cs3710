module decoder_reg
	(
		input rDest_en,
		input [3:0] rDest_in,
		output [15:0] input_out
	)


endmodule

// decoder_reg decode_reg(rDest_en, rDest_in, input_out, regfile_en);